`define DETECT_RISING_EDGE 2'd0
`define DETECT_FALLING_EDGE 2'd1
`define DETECT_BOTH_EDGES 2'd2