`define MY_ENCODER_DECIMAL_DIGIT_WIDTH 4
`define MY_ENCODER_ENCODING_WIDTH 8