`define REG_CTRL_WIDTH 3
`define REG_CTRL_NOP 3'd0
`define REG_CTRL_LD 3'd1
`define REG_CTRL_CLR 3'd2
`define REG_CTRL_INC 3'd3
`define REG_CTRL_DEC 3'd4