`define REG_CTRL_WIDTH 3
`define REG_CTRL_INC 3'b000
`define REG_CTRL_DEC 3'b001
`define REG_CTRL_LD 3'b010
`define REG_CTRL_CLR 3'b011
`define REG_CTRL_NOP 3'b100
