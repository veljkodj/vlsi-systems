`define MY_EDGE_DETECTOR_RISING_EDGE 2'd0
`define MY_EDGE_DETECTOR_FALLING_EDGE 2'd1
`define MY_EDGE_DETECTOR_BOTH_EDGES 2'd2