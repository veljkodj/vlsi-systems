`define MY_ASSOCIATIVE_BUFFER_CTRL_WIDTH 3
`define MY_ASSOCIATIVE_BUFFER_CTRL_NOP 3'd0
`define MY_ASSOCIATIVE_BUFFER_CTRL_CLR 3'd1
`define MY_ASSOCIATIVE_BUFFER_CTRL_LOAD 3'd2
`define MY_ASSOCIATIVE_BUFFER_CTRL_INCR 3'd3